base test 
new line after git git