solarized
colors blue 123
colors red 456
edit after commit
edited in sub1