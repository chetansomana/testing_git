base test 
new line after git add
new line after git commit
